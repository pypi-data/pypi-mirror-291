`ifndef INCLUDED_ZSP_SV_MACROS_SVH
`define INCLUDED_ZSP_SV_MACROS_SVH





`endif /* INCLUDED_ZSP_SV_MACROS_SVH */
